
module multi3();

endmodule

module multi3();

endmodule
