
module multi3();

endmodule

module multi3(p1, p2, result);
	input [2:0] p1;
	input [2:0] p2;

endmodule
